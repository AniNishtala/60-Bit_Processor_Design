module 72_Bit_Processor_Top;

/***************************************************************************/
/************************Wire Instantiate***********************************/
/***************************************************************************/
  wire clk, rst;
  wire Branch_en, Jump_en, immediate_en, read_write_en;
  wire [71:0] Instruction_Fetch;


  /***************************************************************************/
/************************Program Counter Instantiate***********************************/
/***************************************************************************/

  /*
    Program_Counter PC(
      
    );

  */

  
  
endmodule
